`timescale 1ns/1ns
module decode(input [7:0]in,output Q_0,Q_1,Q_2,Q_3,Q_4,Q_5,Q_6,Q_7);
  assign Q_0=in[0];
  assign Q_1=in[1];
  assign Q_2=in[2];
  assign Q_3=in[3];
  assign Q_4=in[4];
  assign Q_5=in[5];
  assign Q_6=in[6];
  assign Q_7=in[7];
endmodule
  
  
  
  
  
  
  

`timescale 1ns/1ns
module Stack(input push,pop,tos,clk,input[7:0] d_in,output[7:0] d_out);
 ...
endmodule
  

`timescale 1ns/1ns
module Memory(input[7:0] writeData,input[4:0] Address,input MemRead,Memwrite,output[7:0] ReadData);
  ...
endmodule  
